module protect(
				

				);
				
				
endmodule