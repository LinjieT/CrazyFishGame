reg[23:0] rand;
  rand = min+{$random}%(max-min+1);